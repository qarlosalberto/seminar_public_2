library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package type_declaration_pkg is
    type t_data is record
        data_0 : std_logic_vector;
        data_1 : std_logic_vector;
    end record t_data;

end package type_declaration_pkg;
